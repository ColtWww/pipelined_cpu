
module vio (
	source,
	probe);	

	output	[0:0]	source;
	input	[0:0]	probe;
endmodule
